module sram #(
    parameter DATA_WIDTH = 64,
    parameter NUM_WORDS  = 1024,
    parameter OUT_REGS   = 0
) (
    input  logic                         clk_i,
    input  logic                         rst_ni,
    input  logic                         req_i,
    input  logic                         we_i,
    input  logic [$clog2(NUM_WORDS)-1:0] addr_i,
    input  logic [       DATA_WIDTH-1:0] wdata_i,
    input  logic [ (DATA_WIDTH+7)/8-1:0] be_i,
    output logic [       DATA_WIDTH-1:0] rdata_o
);

  localparam DATA_WIDTH_ALIGNED = ((DATA_WIDTH + 63) / 64) * 64;
  localparam BE_WIDTH_ALIGNED = (((DATA_WIDTH + 7) / 8 + 7) / 8) * 8;

  logic [DATA_WIDTH_ALIGNED-1:0] wdata_aligned;
  logic [  BE_WIDTH_ALIGNED-1:0] be_aligned;
  logic [DATA_WIDTH_ALIGNED-1:0] rdata_aligned;

  always_comb begin : p_align
    wdata_aligned                    = '0;
    be_aligned                       = '0;
    wdata_aligned[DATA_WIDTH-1:0]    = wdata_i;
    be_aligned[BE_WIDTH_ALIGNED-1:0] = be_i;

    rdata_o                          = rdata_aligned[DATA_WIDTH-1:0];
  end

  genvar k;
  generate
    for (k = 0; k < (DATA_WIDTH + 63) / 64; k++) begin

      SyncSpRamBeNx64 #(
          .ADDR_WIDTH($clog2(NUM_WORDS)),
          .DATA_DEPTH(NUM_WORDS),
          .OUT_REGS  (0),
          .SIM_INIT  (2)
      ) i_ram (
          .Clk_CI   (clk_i),
          .Rst_RBI  (rst_ni),
          .CSel_SI  (req_i),
          .WrEn_SI  (we_i),
          .BEn_SI   (be_aligned[k*8+:8]),
          .WrData_DI(wdata_aligned[k*64+:64]),
          .Addr_DI  (addr_i),
          .RdData_DO(rdata_aligned[k*64+:64])
      );
    end
  endgenerate

endmodule : sram
